
//=====================================================================
//
// Description:
//  The files to include all the macro defines
//
// ====================================================================


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////// ISA relevant macro
//
`define QPDAC_INSTR_SIZE 32
`define QPDAC_ITCM_WIDTH 32
//////////////////////////test//////////////////
//`define QPDAC_PC_SIZE 11
/////////////////////////test///////////////////
`define QPDAC_PC_SIZE 14


`define QPDAC_ADDR_SIZE 14
`define QPDAC_REPEAT_LEN 28

`define QPDAC_DATA_WIDTH  32                           

`define QPDAC_QXLEN 31

`define QPDAC_REPEAT_STACK_DEPTH 8

 `define QPDAC_DECINFO_GRP_WIDTH    2
  `define QPDAC_DECINFO_GRP_ALU      `QPDAC_DECINFO_GRP_WIDTH'd1
  `define QPDAC_DECINFO_GRP_BJP      `QPDAC_DECINFO_GRP_WIDTH'd2
  `define QPDAC_DECINFO_GRP_QIU      `QPDAC_DECINFO_GRP_WIDTH'd3
  
      `define QPDAC_DECINFO_GRP_LSB  0
      `define QPDAC_DECINFO_GRP_MSB  (`QPDAC_DECINFO_GRP_LSB+`QPDAC_DECINFO_GRP_WIDTH-1)
  `define QPDAC_DECINFO_GRP          `QPDAC_DECINFO_GRP_MSB:`QPDAC_DECINFO_GRP_LSB
  
  `define QPDAC_DECINFO_SUBDECINFO_LSB    (`QPDAC_DECINFO_GRP_MSB+1)

  
  
// ALU group
      `define QPDAC_DECINFO_ALU_IMM_LSB    `QPDAC_DECINFO_SUBDECINFO_LSB
      `define QPDAC_DECINFO_ALU_IMM_MSB    (`QPDAC_DECINFO_ALU_IMM_LSB+`QPDAC_REPEAT_LEN-1)
  `define QPDAC_DECINFO_ALU_IMM    `QPDAC_DECINFO_ALU_IMM_MSB :`QPDAC_DECINFO_ALU_IMM_LSB 
       `define QPDAC_DECINFO_ALU_WIDTH    (`QPDAC_DECINFO_ALU_IMM_MSB+1)


  // Bxx group
      `define QPDAC_DECINFO_BJP_BPRDT_LSB `QPDAC_DECINFO_SUBDECINFO_LSB
      `define QPDAC_DECINFO_BJP_BPRDT_MSB (`QPDAC_DECINFO_BJP_BPRDT_LSB+1-1)
  `define QPDAC_DECINFO_BJP_BPRDT  `QPDAC_DECINFO_BJP_BPRDT_MSB:`QPDAC_DECINFO_BJP_BPRDT_LSB
      `define QPDAC_DECINFO_BJP_CMP_LSB (`QPDAC_DECINFO_BJP_BPRDT_MSB+1)
      `define QPDAC_DECINFO_BJP_CMP_MSB (`QPDAC_DECINFO_BJP_CMP_LSB+1-1)
  `define QPDAC_DECINFO_BJP_CMP    `QPDAC_DECINFO_BJP_CMP_MSB  :`QPDAC_DECINFO_BJP_CMP_LSB  
      `define QPDAC_DECINFO_BJP_REPEAT_LSB (`QPDAC_DECINFO_BJP_CMP_MSB+1)
      `define QPDAC_DECINFO_BJP_REPEAT_MSB (`QPDAC_DECINFO_BJP_REPEAT_LSB+1-1)
  `define QPDAC_DECINFO_BJP_REPEAT    `QPDAC_DECINFO_BJP_REPEAT_MSB  :`QPDAC_DECINFO_BJP_REPEAT_LSB  
      `define QPDAC_DECINFO_BJP_GOTO_LSB (`QPDAC_DECINFO_BJP_REPEAT_MSB+1)
      `define QPDAC_DECINFO_BJP_GOTO_MSB (`QPDAC_DECINFO_BJP_GOTO_LSB+1-1)
  `define QPDAC_DECINFO_BJP_GOTO    `QPDAC_DECINFO_BJP_GOTO_MSB  :`QPDAC_DECINFO_BJP_GOTO_LSB  
      `define QPDAC_DECINFO_BJP_IMM_LSB (`QPDAC_DECINFO_BJP_GOTO_MSB+1)
      `define QPDAC_DECINFO_BJP_IMM_MSB (`QPDAC_DECINFO_BJP_IMM_LSB+`QPDAC_ADDR_SIZE-1)
  `define QPDAC_DECINFO_BJP_IMM    `QPDAC_DECINFO_BJP_IMM_MSB  :`QPDAC_DECINFO_BJP_IMM_LSB  
  
`define QPDAC_DECINFO_BJP_WIDTH  (`QPDAC_DECINFO_BJP_IMM_MSB+1)

  //Quantum Instruction group
      `define QPDAC_DECINFO_QIU_PARA_LSB `QPDAC_DECINFO_SUBDECINFO_LSB
      `define QPDAC_DECINFO_QIU_PARA_MSB (`QPDAC_DECINFO_QIU_PARA_LSB + `QPDAC_QXLEN - 1)
    `define QPDAC_DECINFO_QIU_PARA  `QPDAC_DECINFO_QIU_PARA_MSB : `QPDAC_DECINFO_QIU_PARA_LSB
    
`define QPDAC_DECINFO_QIU_WIDTH  (`QPDAC_DECINFO_QIU_PARA_MSB+1)

`define QPDAC_DECINFO_WIDTH  `QPDAC_DECINFO_QIU_WIDTH



`define FEEDBACK 1'b1

`define CPU_WF_ADDR_SIZE  17
`define CPU_WF_DURATION_SIZE 10
`define CPU_WF_MODE_SIZE 4
`define CPU_WF_TRIGGER_SIZE 1
`define CPU_WF_TYPE_SIZE 2
`define CPU_WF_SEL_SIZE 1


`define WF_ADDR_SIZE 10
`define WF_AMP_SIZE 17
`define WF_DURATION_SIZE 10
`define WF_MODE_SIZE 3
`define WF_SEL_SIZE 1
`define WF_TRIGGER_SIZE 1
`define WF_TYPE_SIZE 2
`define WF_INSTR_SIZE  (`WF_AMP_SIZE + `WF_DURATION_SIZE + `WF_MODE_SIZE +`WF_TRIGGER_SIZE + `WF_TRIGGER_SIZE + `WF_TYPE_SIZE)


`define WF_INSTR_BUFF_DEPTH 32
`define WF_WVFORM_FIFO_DEPTH 16

`define WF_SEL_SIZE 1
`define WF_DEFMODE_SIZE 1
`define WF_SET_MODE_TYPE_SIZE 2

`define WF_TYPE_IN_MODE  (`WF_DEFMODE_SIZE + `WF_SET_MODE_TYPE_SIZE - 1) :`WF_DEFMODE_SIZE
`define WF_DEFMODE_IN_MODE (`WF_DEFMODE_SIZE - 1) : 0
`define WF_SEL_IN_MODE (`WF_SEL_SIZE - 1) : 0

`define WF_INSTR_EXU_ODATA_SIZE (`WF_INSTR_EXU_ODATA_TYPE_SEL_SIZE + `WF_MODE_SIZE + `WF_AMP_SIZE)                              //////{type_is_setmode , type_is_wait, mode, amp}
`define WF_INSTR_EXU_ODATA_TYPE_SEL_SIZE 2                                                               /////type_is_setmode , type_is_wait

`define WF_DEF_LENGTH_SIZE 12




    `define CPU_WF_DATA_LSB 0
    `define CPU_WF_DATA_MSB (`CPU_WF_DATA_LSB + `CPU_WF_ADDR_SIZE - 1)
`define CPU_WF_DATA `CPU_WF_DATA_MSB :  `CPU_WF_DATA_LSB
 
    `define CPU_WF_DURATION_LSB (`CPU_WF_DATA_MSB + 1)
    `define CPU_WF_DURATION_MSB (`CPU_WF_DURATION_LSB + `CPU_WF_DURATION_SIZE - 1)
`define CPU_WF_DURATION `CPU_WF_DURATION_MSB :  `CPU_WF_DURATION_LSB

    `define CPU_WF_MODE_LSB (`CPU_WF_DURATION_MSB + 1)
    `define CPU_WF_MODE_MSB (`CPU_WF_MODE_LSB + `CPU_WF_MODE_SIZE - 1)
`define CPU_WF_MODE `CPU_WF_MODE_MSB :  `CPU_WF_MODE_LSB

    `define CPU_WF_TRIGGER_LSB (`CPU_WF_MODE_MSB + 1)
    `define CPU_WF_TRIGGER_MSB (`CPU_WF_TRIGGER_LSB + `CPU_WF_TRIGGER_SIZE - 1)
`define CPU_WF_TRIGGER `CPU_WF_TRIGGER_MSB :  `CPU_WF_TRIGGER_LSB


    `define CPU_WF_TYPE_LSB (`CPU_WF_TRIGGER_MSB + 1)
    `define CPU_WF_TYPE_MSB (`CPU_WF_TYPE_LSB + `CPU_WF_TYPE_SIZE - 1)
`define CPU_WF_TYPE `CPU_WF_TYPE_MSB :  `CPU_WF_TYPE_LSB

    `define CPU_WF_SEL_LSB `CPU_WF_MODE_LSB
    `define CPU_WF_SEL_MSB (`CPU_WF_MODE_LSB + `CPU_WF_SEL_SIZE - 1)
`define CPU_WF_SEL `CPU_WF_SEL_MSB : `CPU_WF_SEL_LSB    




    `define WF_DATA_LSB 0
    `define WF_DATA_MSB (`WF_DATA_LSB + `WF_ADDR_SIZE - 1)
`define WF_DATA `WF_DATA_MSB :  `WF_DATA_LSB
 
    `define WF_DURATION_LSB (`WF_DATA_MSB + 1)
    `define WF_DURATION_MSB (`WF_DURATION_LSB + `WF_DURATION_SIZE - 1)
`define WF_DURATION `WF_DURATION_MSB :  `WF_DURATION_LSB

    `define WF_MODE_LSB (`WF_DURATION_MSB + 1)
    `define WF_MODE_MSB (`WF_MODE_LSB + `WF_MODE_SIZE - 1)
`define WF_MODE `WF_MODE_MSB :  `WF_MODE_LSB

    `define WF_TRIGGER_LSB (`WF_MODE_MSB + 1)
    `define WF_TRIGGER_MSB (`WF_TRIGGER_LSB + `WF_TRIGGER_SIZE - 1)
`define WF_TRIGGER `WF_TRIGGER_MSB :  `WF_TRIGGER_LSB


    `define WF_TYPE_LSB (`WF_TRIGGER_MSB + 1)
    `define WF_TYPE_MSB (`WF_TYPE_LSB + `WF_TYPE_SIZE - 1)
`define WF_TYPE `WF_TYPE_MSB :  `WF_TYPE_LSB




    `define WF_INSTR_EXU_ODATA_DATA_LSB 0
    `define WF_INSTR_EXU_ODATA_DATA_MSB  (`WF_INSTR_EXU_ODATA_DATA_LSB  + `WF_AMP_SIZE - 1)
`define WF_INSTR_EXU_ODATA_DATA `WF_INSTR_EXU_ODATA_DATA_MSB :  `WF_INSTR_EXU_ODATA_DATA_LSB
 
    `define WF_INSTR_EXU_ODATA_MODE_LSB (`WF_INSTR_EXU_ODATA_DATA_MSB + 1)
    `define WF_INSTR_EXU_ODATA_MODE_MSB (`WF_INSTR_EXU_ODATA_MODE_LSB + `WF_MODE_SIZE - 1)
`define WF_INSTR_EXU_ODATA_MODE `WF_INSTR_EXU_ODATA_MODE_MSB :  `WF_INSTR_EXU_ODATA_MODE_LSB

    `define WF_INSTR_EXU_ODATA_TYPE_SEL_LSB (`WF_INSTR_EXU_ODATA_MODE_MSB + 1)
    `define WF_INSTR_EXU_ODATA_TYPE_SEL_MSB (`WF_INSTR_EXU_ODATA_TYPE_SEL_LSB + `WF_INSTR_EXU_ODATA_TYPE_SEL_SIZE - 1)
`define WF_INSTR_EXU_ODATA_TYPE_SEL `WF_INSTR_EXU_ODATA_TYPE_SEL_MSB :  `WF_INSTR_EXU_ODATA_TYPE_SEL_LSB


`define INS_MEM_BROM_NUM 1
`define WF_MEM_HROM_NUM 1
`define LENGTH_MEM_HROM_NUM 2
`define DEF_MEM_HROM_NUM 3

`define BROM_DIR "E:/gitlab/distribution-quantum-architecture/BROM"
`define HROM_DIR "E:/gitlab/distribution-quantum-architecture/HROM"
`define ROM_FILE_TYPE ".txt"
//////////////
`define DATA_WIDTH 64

/////////////////DATA WIDTH IN PC INSTRUCTION
`define INS_TYPE_WIDTH 8
`define TASK_ID_WIDTH 8
`define TASK_NUMBER_WIDTH 8
`define CHANNEL_NUMBER_WIDTH 8

`define DAC_CHANNEL_MASK_WIDTH 8
`define DAC_UNDEFINE_WIDTH 16
`define DAC_TASK_TYPE_WIDTH 8

///////////////TASK ADDR WRITE MODULE
`define DAC_TASKADDR_WIDTH 64
`define DAC_TASKADDR_ADDR_WIDTH 4

//////////////WAVEFORM WRITE MODULE
`define DAC_TASK_WF_DATA_WIDTH 512
`define DAC_TASK_WF_DATAADDR_WIDTH 16
`define DAC_TASK_WF_INSADDR_WIDTH 16

`define DAC_WFWR_CHANNEL_MASK_INS_WIDTH 32
`define DAC_WFWR_CHANNEL_MASK_WIDTH 4
`define DAC_WFWR_WF_LENGTH_WIDTH 16
`define DAC_WFWR_CYCLE_NUM_WIDTH 16


//////////////TASK CORE TOP
`define DAC_TASKCORE_TASK_MUMBER_WIDTH 4

/////////////DAC CONF MODULE
`define DAC_TRIGGER_LENGTH 5'd5
`define DAC_TRIGGER_CYCLE  8'd50
`define DAC_SYNC_LENGTH  5'd10

////////////waveform_play module
`define DAC_WF_ADDR_WIDTH 12
`define DAC_WF_VALIDDATA_WIDTH 384
`define DAC_WF_VALIDDATA_TO_DAC_WIDTH 128


    `define INS_TYPE_LSB 0
    `define INS_TYPE_MSB (`INS_TYPE_LSB + `INS_TYPE_WIDTH - 1)
`define INS_TYPE `INS_TYPE_MSB :  `INS_TYPE_LSB
 
    `define TASK_ID_LSB (`INS_TYPE_MSB + 1)
    `define TASK_ID_MSB (`TASK_ID_LSB + `TASK_ID_WIDTH - 1)
`define TASK_ID `TASK_ID_MSB :  `TASK_ID_LSB

    `define DAC_CHANNEL_MASK_LSB (`TASK_ID_MSB + 1)
    `define DAC_CHANNEL_MASK_MSB (`DAC_CHANNEL_MASK_LSB + `DAC_CHANNEL_MASK_WIDTH - 1)
`define DAC_CHANNEL_MASK `DAC_CHANNEL_MASK_MSB :  `DAC_CHANNEL_MASK_LSB

    `define DAC_UNDEFINE_LSB (`DAC_CHANNEL_MASK_MSB + 1)
    `define DAC_UNDEFINE_MSB (`DAC_UNDEFINE_LSB + `DAC_UNDEFINE_WIDTH - 1)
`define DAC_UNDEFINE `DAC_UNDEFINE_MSB :  `DAC_UNDEFINE_LSB

    `define TASK_NUMBER_LSB (`DAC_UNDEFINE_MSB + 1)
    `define TASK_NUMBER_MSB (`TASK_NUMBER_LSB + `TASK_NUMBER_WIDTH - 1)
`define TASK_NUMBER `TASK_NUMBER_MSB :  `TASK_NUMBER_LSB

    `define DAC_TASK_TYPE_LSB (`TASK_NUMBER_MSB + 1)
    `define DAC_TASK_TYPE_MSB (`DAC_TASK_TYPE_LSB + `DAC_TASK_TYPE_WIDTH - 1)
`define DAC_TASK_TYPE `DAC_TASK_TYPE_MSB :  `DAC_TASK_TYPE_LSB

    `define CHANNEL_NUMBER_LSB (`DAC_TASK_TYPE_MSB + 1)
    `define CHANNEL_NUMBER_MSB (`CHANNEL_NUMBER_LSB + `CHANNEL_NUMBER_WIDTH - 1)
`define CHANNEL_NUMBER `CHANNEL_NUMBER_MSB :  `CHANNEL_NUMBER_LSB

//////////////DAC WF WR MODULE
    `define DAC_WFWR_CHANNEL_MASK_LSB 0
    `define DAC_WFWR_CHANNEL_MASK_MSB (`DAC_WFWR_CHANNEL_MASK_LSB + `DAC_WFWR_CHANNEL_MASK_INS_WIDTH - 1)
`define DAC_WFWR_CHANNEL_MASK `DAC_WFWR_CHANNEL_MASK_MSB :  `DAC_WFWR_CHANNEL_MASK_LSB
 
    `define DAC_WFWR_WF_LENGTH_LSB (`DAC_WFWR_CHANNEL_MASK_MSB + 1)
    `define DAC_WFWR_WF_LENGTH_MSB (`DAC_WFWR_WF_LENGTH_LSB + `DAC_TASK_WF_DATAADDR_WIDTH - 1)
`define DAC_WFWR_WF_LENGTH `DAC_WFWR_WF_LENGTH_MSB :  `DAC_WFWR_WF_LENGTH_LSB

    `define DAC_WFWR_INS_LENGTH_LSB (`DAC_WFWR_WF_LENGTH_MSB + 1)
    `define DAC_WFWR_INS_LENGTH_MSB (`DAC_WFWR_INS_LENGTH_LSB + `DAC_TASK_WF_INSADDR_WIDTH - 1)
`define DAC_WFWR_INS_LENGTH `DAC_WFWR_INS_LENGTH_MSB :  `DAC_WFWR_INS_LENGTH_LSB

////////////////////////////
`define ADDA_WF_ADDR_WIDTH 9
`define ADDA_WF_DATA_WIDTH 512 //8
`define ADDA_WF_VALID_DATA_WIDTH 384///16

`define ADDA_QUBIT_NUMBER_PER_CHANNEL 6///2
`define ADDA_CHANNEL_NUMBER 4
`define ADDA_QUBIT_NUMBER (`ADDA_CHANNEL_NUMBER * `ADDA_QUBIT_NUMBER_PER_CHANNEL)

`define ADDA_CONFIG_NUMBER_WIDTH 8
`define ADDA_CONFIG_CHANNEL_NUMBER_WIDTH 8

`define ADDA_CONFIGADDR_WIDTH 64
`define ADDA_CONFIGADDR_ADDR_WIDTH 4

`define ADDA_TASKADDR_ADDR_WIDTH 4
`define ADDA_TASKADDR_WIDTH 64

`define ADDA_CYCLE_NUM_WIDTH 16
`define ADDA_TIMING_INS_ADDR_WIDTH 4
`define ADDA_TIMING_INS_DATA_WIDTH 32
`define ADDA_MEASURE_TIMES_WIDTH 8

`define ADDA_TIMEING_COUNTER_WIDTH 16

`define ADDA_WF_VALIDDATA_TO_ADDA_WIDTH 128
`define ADDA_SAMPLE_NUMBER 32
`define ADDA_SAMPLE_WIDTH 12




`define ADDA_FACTOR_DATA_WIDTH 512
`define ADDA_FACTOR_VALID_DATA_WIDTH 480           
`define ADDA_FACTOR_ADDR_WIDTH 9

`define ADDA_ORIGIN_DATA_WIDTH 480///32
`define ADDA_ORIGIN_DATA_ADDR_WIDTH 11

`define ADDA_IQ_DATA_WIDTH 32//8
`define ADDA_IQ_DATA_ADDR_WIDTH 4

`define ADDA_WORK_MODE_WIDTH 2

`define ADDA_TASK_WB_DATA_LENGTH_WIDTH 32
`define ADDA_SINGLE_WB_DATA_LENGTH_WIDTH 16
`define ADDA_CHANNEL_WB_DATA_LENGTH_WIDTH 24

`define ADDA_USED_FACTOR_ADDR_WIDTH 4
`define ADDA_SIMPLE_ADDR_WIDTH 12




`define DDR_ADDR_WIDTH  28


`define ORIGIN_DATA_MEM_MAX_ADDR 1600

`define FACTOR_DATA_MEM_MAX_ADDR 320

`define IQ_DATA_MEM_MAX_ADDR 16

`define DDR_DATA_WIDTH 512

`define BUFFER_DATA_LENGTH_WIDTH 12

`define TASKCORE_NUM 1
`define DDR_NUM 2
`define ADDA_CHANNEL_NUMBER_PER_DDR  (`ADDA_CHANNEL_NUMBER / `DDR_NUM)

`define AURORA_DATA_WIDTH 64
`define VPX_NUM_WIDTH 8